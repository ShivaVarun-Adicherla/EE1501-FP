module top_module();
initial begin
  $display("Hello World");
endmodule
