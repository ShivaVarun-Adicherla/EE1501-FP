module time_to 
